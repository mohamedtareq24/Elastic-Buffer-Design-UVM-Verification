`define DATA_WIDTH 20
`define FIFO_DEPTH 