package eb_common_pkg;
  // Global SKP ordered set constants (K28.1 & K28.1 with alternating disparity)
  parameter bit [19:0] USB_SKP_VAL_1 = {10'b1100000110, 10'b0011111001};
  parameter bit [19:0] USB_SKP_VAL_2 = {10'b0011111001, 10'b1100000110};
endpackage : eb_common_pkg
