package rd_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "rd_item.sv"
  `include "rd_mon_tr.sv"
// `include "rd_sequencer.sv"
//`include "rd_driver.sv"
  `include "rd_monitor.sv"
  `include "rd_agent.sv"
//`include "rd_base_seq.sv"

endpackage : rd_pkg
